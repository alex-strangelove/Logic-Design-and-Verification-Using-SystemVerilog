`timescale 1ns/1ps

module fourBitTest(output logic a, b, c, d);
endmodule: fourBitTest