`timescale 1ns/1ns

module fourBitTest
(
    input logic a, b, c, d
);
endmodule: fourBitTest